fbgjnk
